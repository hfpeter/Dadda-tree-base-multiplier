
module dadda_tree (b_3bit,p,S);

input [11:0] p[0:6];
output [21:0] S; 

input [2:0] b_3bit [0:6];
wire [2:0] b_3bit [0:6];

wire [11:0] p[0:6];
wire [5 :0]  q0 ; 
wire [13 :0] q1 ; 
wire [9 :0] q2 ; 
wire [17:0] q3 ; 
wire [20:0] q4 ; 
wire [23:0] q5 ; 
wire [5 :0] c0 ;
wire [13  :0] c1 ; 
wire [9:0] c2 ; 
wire [17:0] c3 ; 
wire [20:0] c4 ; 
wire [23:0] c5 ; 
wire ns0; 
wire ns1; 
wire ns2;
wire ns3;
wire ns4 ; 
wire ns5; 
wire s0; 
wire s1; 
wire s2;
wire s3;
wire s4 ; 
wire s5; 
assign s0=b_3bit[0][2];
assign s1=b_3bit[1][2];
assign s2=b_3bit[2][2];
assign s3=b_3bit[3][2];
assign s4=b_3bit[4][2];
assign s5=b_3bit[5][2];

assign ns0=~b_3bit[0][2]; 
assign ns1=~b_3bit[1][2]; 
assign ns2=~b_3bit[2][2]; 
assign ns3=~b_3bit[3][2]; 
assign ns4=~b_3bit[4][2]; 
assign ns5=~b_3bit[5][2]; 
HA	F0 (p[0][10],p[1][8],q0[0]	,c0[0]	);
HA	F1 (p[0][11],p[1][9],q0[1]	,c0[1]	);
FA	F2 (s0	,p[1][10],p[2][8],q0[2]	,c0[2]	);
FA	F3 (s0	,p[1][11],p[2][9],q0[3]	,c0[3]	);
FA	F4 (ns0	,ns1	 ,p[2][10],q0[4]	,c0[4]	);
HA	F5 (1'b1	,p[2][11],q0[5]	,c0[5]	);

HA	F7 (p[0][6]	,p[1][4] ,q1[0 ]	,c1[0 ]	);	
HA	F8 (p[0][7]	,p[1][5] ,q1[1 ]	,c1[1 ]	);	
FA	F9 (p[0][8]	,p[1][6] ,p[2][4]	,q1[2 ]	,c1[2 ]	);HA	F62(p[3][2],p[4][0],q2[0]	,c2[0]);
FA	F10(p[0][9]	,p[1][7] ,p[2][5]	,q1[3 ]	,c1[3 ]	);HA	F63(p[3][3],p[4][1],q2[1]	,c2[1]);
FA	F11(q0[0]	,p[2][6] ,p[3][4],q1[4 ]	,c1[4 ]	);	FA	F64(p[4][2],p[5][0],	s5,q2[2]	,c2[2]);
FA	F12(c0[0]	,q0[1]	 ,p[2][7],q1[5 ]	,c1[5 ]	);	FA	F65(p[3][5],p[4][3],	p[5][1],q2[3]	,c2[3]);
FA	F13(c0[1]	,q0[2]	 ,p[3][6],q1[6 ]	,c1[6 ]	);	FA	F66(p[4][4],p[5][2],	p[6][0],q2[4]	,c2[4]);
FA	F14(c0[2]	,q0[3]	 ,p[3][7],q1[7 ]	,c1[7 ]	);	FA	F67(p[4][5],p[5][3],	p[6][1],q2[5]	,c2[5]);
FA	F15(c0[3]	,q0[4]	 ,p[3][8],q1[8 ]	,c1[8 ]	);	FA	F68(p[4][6],p[5][4],	p[6][2],q2[6]	,c2[6]);
FA	F16(c0[4]	,q0[5]	 ,p[3][9],q1[9 ]	,c1[9 ]	);	FA	F69(p[4][7],p[5][5],	p[6][3],q2[7]	,c2[7]);
FA	F17(c0[5]	,ns2	 ,p[3][10],q1[10]	,c1[10]	);	FA	F70(p[4][8],p[5][6],	p[6][4],q2[8]	,c2[8]);
FA	F18(1'b1	,p[3][11],p[4][9],q1[11]	,c1[11]	);      HA	F71(p[5][7],p[6][5],q2[9]	,c2[9]);
FA	F19(ns3	,p[4][10],p[5][8],q1[12]	,c1[12]	);
HA	F20(1'b1	,p[4][11],q1[13]	,c1[13]	);

HA	F22(p[0][4]	,p[1][2] , q3[0 ]	,c3[0 ]	);
HA	F23(p[0][5]	,p[1][3] , q3[1 ]	,c3[1 ]	);
FA	F24(q1[0]	,p[2][2] ,p[3][0],q3[2 ]	,c3[2 ]	);
FA	F25(c1[0 ]	,q1[1]	 ,p[2][3],q3[3 ]	,c3[3 ]	);
FA	F26(c1[1 ]	,q1[2]	 ,q2[0],q3[4 ]	,c3[4 ]	);
FA	F27(c1[2 ]	,c2[0]	 ,q1[3],q3[5 ]	,c3[5 ]	);
FA	F28(c1[3 ]	,c2[1]	 ,q1[4],q3[6 ]	,c3[6 ]	);
FA	F29(c1[4 ]	,c2[2]	 ,q1[5],q3[7 ]	,c3[7 ]	);
FA	F30(c1[5 ]	,c2[3]	 ,q1[6],q3[8 ]	,c3[8 ]	);
FA	F31(c1[6 ]	,c2[4]	 ,q1[7],q3[9 ]	,c3[9 ]	);
FA	F32(c1[7 ]	,c2[5]	 ,q1[8],q3[10]	,c3[10]	);
FA	F33(c1[8 ]	,c2[6]	 ,q1[9],q3[11]	,c3[11]	);
FA	F34(c1[9 ]	,c2[7]	 ,q1[10],q3[12]	,c3[12]	);
FA	F35(c1[10]	,c2[8]	 ,q1[11],q3[13]	,c3[13]	);
FA	F36(c1[11]	,c2[9]	 ,q1[12],q3[14]	,c3[14]	);
FA	F37(c1[12]	,q1[13]	 ,p[5][9],q3[15]	,c3[15]	);
FA	F38(c1[13]	,ns4	 ,p[5][10],q3[16]	,c3[16]	);
HA	F39(1'b1	,p[5][11],q3[17]	,c3[17]	);

HA	F41(p[0][2]	,p[1][0],q4[0 ]	,c4[0 ]	);
HA	F42(p[0][3]	,p[1][1],q4[1 ]	,c4[1 ]	);
FA	F43(q3[0]	,p[2][0] ,s2,q4[2 ]	,c4[2 ]	);
FA	F44(c3[0 ]	,q3[1 ]	 ,p[2][1],q4[3 ]	,c4[3 ]	);
FA	F45(c3[1 ]	,q3[2 ]	 ,s3,q4[4 ]	,c4[4 ]	);
FA	F46(c3[2 ]	,q3[3 ]	 ,p[3][1],q4[5 ]	,c4[5 ]	);
FA	F47(c3[3 ]	,q3[4 ]	 ,s4   ,q4[6 ]	,c4[6 ]	);
FA	F48(c3[4 ]	,q3[5 ]	 ,q2[1],q4[7 ]	,c4[7 ]	);
FA	F49(c3[5 ]	,q3[6 ]	 ,q2[2],q4[8 ]	,c4[8 ]	);
FA	F50(c3[6 ]	,q3[7 ]	 ,q2[3],q4[9 ]	,c4[9 ]	);
FA	F51(c3[7 ]	,q3[8 ]	 ,q2[4],q4[10]	,c4[10]	);
FA	F52(c3[8 ]	,q3[9 ]	 ,q2[5],q4[11]	,c4[11]	);
FA	F53(c3[9 ]	,q3[10]	 ,q2[6],q4[12]	,c4[12]	);
FA	F54(c3[10]	,q3[11]	 ,q2[7],q4[13]	,c4[13]	);
FA	F55(c3[11]	,q3[12]	 ,q2[8],q4[14]	,c4[14]	);
FA	F56(c3[12]	,q3[13]	 ,q2[9],q4[15]	,c4[15]	);
FA	F57(c3[13]	,q3[14]	 ,p[6][6],q4[16]	,c4[16]	);
FA	F58(c3[14]	,q3[15]	 ,p[6][7],q4[17]	,c4[17]	);
FA	F59(c3[15]	,q3[16]	 ,p[6][8],q4[18]	,c4[18]	);
FA	F60(c3[16]	,q3[17]	 ,p[6][9],q4[19]	,c4[19]	);
FA	F61(c3[17]	,ns5	 ,p[6][10],q4[20]	,c4[20]	);

HA AF0(p[0][0	] , s0,                  q5[0],c5[0]);
FA	A161n	( p[0][1	] ,	1'b0 ,	c5[0] ,  q5[1],c5[1]);
FA	A161m	( q4[0	] ,	s1 ,	c5[1] ,  q5[2],c5[2]);

    genvar i;
    generate
    for (i = 0; i <=19; i = i + 1) begin
    FA	A161b	( c4[i] ,q4[i+1] ,c5[i+2] , q5[i+3],c5[i+3]);
    end
    endgenerate
HA AF1(c4[20] , c5[22],                  q5[23],c5[23]);
 assign S[21:0]=q5[21:0];
endmodule

